 Hi this is Nagaraju sadanandan file
