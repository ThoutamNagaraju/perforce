 Hi this is Nagaraju sadanandan file-edited1
