 Hi this is Nagaraju sadanandan file-edited1
 Hi this is Nagaraju sadanandan file-edited2
